`timescale 1ns / 1ps

module clock_consumer_sv (
    // Master signals
    input logic clk

);
endmodule
