entity clock_consumer_v2 is
	port (
		clk 		: in bit
	);
end clock_consumer_v2;

architecture arch_consume of clock_consumer_v2 is
begin

end arch_consume;

