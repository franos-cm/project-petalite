entity clock_consumer_vhd is
	port (
		clk 		: in bit
	);
end clock_consumer_vhd;

architecture arch_consume of clock_consumer_vhd is
begin

end arch_consume;

